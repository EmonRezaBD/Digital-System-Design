CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 108 262 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44092.5 0
0
13 Logic Switch~
5 110 205 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44092.5 0
0
5 4049~
219 644 217 0 2 22
0 6 5
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3124 0 0
2
44092.5 0
0
14 Logic Display~
6 871 341 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
44092.5 0
0
14 Logic Display~
6 865 188 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
44092.5 0
0
10 2-In NAND~
219 361 367 0 3 22
0 3 2 4
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5572 0 0
2
44092.5 0
0
9 2-In AND~
219 359 222 0 3 22
0 3 2 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8901 0 0
2
44092.5 0
0
7
0 2 2 0 0 8192 0 0 6 6 0 3
213 262
213 376
337 376
0 1 3 0 0 8192 0 0 6 7 0 3
178 205
178 358
337 358
3 1 4 0 0 4224 0 6 4 0 0 3
388 367
871 367
871 359
2 1 5 0 0 4224 0 3 5 0 0 3
665 217
865 217
865 206
3 1 6 0 0 4224 0 7 3 0 0 4
380 222
621 222
621 217
629 217
1 2 2 0 0 4224 0 1 7 0 0 4
120 262
327 262
327 231
335 231
1 1 3 0 0 4224 0 2 7 0 0 4
122 205
327 205
327 213
335 213
13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
816 459 901 483
826 467 890 483
8 switches
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
933 437 1122 461
943 445 1111 461
21 input, then connect n
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
816 436 941 460
826 444 930 460
13 if there is n
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
948 415 1097 439
958 423 1086 439
16 input NAND gates
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
809 414 958 438
819 422 947 438
16 *Same for 3 or 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
911 328 1092 352
921 336 1081 352
20 Using NAND Gate Chip
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
893 181 1050 205
903 189 1039 205
17 Using Basic Gates
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
443 426 576 450
453 434 565 450
14 Fig: NAND Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
535 332 596 356
545 340 585 356
5 (AB)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
743 183 804 207
753 191 793 207
5 (AB)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
461 179 498 203
471 187 487 203
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
93 273 122 297
103 281 111 297
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
94 128 123 152
104 136 112 152
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
