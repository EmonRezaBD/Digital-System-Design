CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 60 30 100 10
176 80 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 423 103 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
44080.8 0
0
13 Logic Switch~
5 281 106 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7876 0 0
2
44080.8 0
0
13 Logic Switch~
5 165 108 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6369 0 0
2
44080.8 0
0
14 Logic Display~
6 1105 521 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9172 0 0
2
44080.8 0
0
8 3-In OR~
219 967 712 0 4 22
0 5 4 3 2
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
7100 0 0
2
44080.8 0
0
9 2-In AND~
219 722 805 0 3 22
0 7 6 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3820 0 0
2
44080.8 0
0
9 2-In AND~
219 723 712 0 3 22
0 7 8 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
7678 0 0
2
44080.8 0
0
9 2-In AND~
219 722 613 0 3 22
0 6 8 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
961 0 0
2
44080.8 0
0
8 2-In OR~
219 1026 372 0 3 22
0 11 10 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3178 0 0
2
44080.8 0
0
9 2-In AND~
219 965 468 0 3 22
0 13 12 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3409 0 0
2
44080.8 0
0
9 2-In AND~
219 946 265 0 3 22
0 14 7 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3951 0 0
2
44080.8 0
0
14 Logic Display~
6 1097 356 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8885 0 0
2
44080.8 0
0
8 2-In OR~
219 832 459 0 3 22
0 16 15 13
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3780 0 0
2
44080.8 0
0
9 2-In AND~
219 724 520 0 3 22
0 6 8 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9265 0 0
2
44080.8 0
0
9 2-In AND~
219 723 422 0 3 22
0 18 17 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9442 0 0
2
44080.8 0
0
8 2-In OR~
219 830 256 0 3 22
0 20 19 14
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9424 0 0
2
44080.8 0
0
9 2-In AND~
219 719 306 0 3 22
0 6 17 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9968 0 0
2
44080.8 0
0
9 2-In AND~
219 714 216 0 3 22
0 18 8 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9281 0 0
2
44080.8 0
0
9 Inverter~
13 491 134 0 2 22
0 8 17
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
8464 0 0
2
44080.8 0
0
9 Inverter~
13 342 136 0 2 22
0 6 18
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7168 0 0
2
44080.8 0
0
9 Inverter~
13 199 141 0 2 22
0 12 7
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3171 0 0
2
44080.8 0
0
32
4 1 2 0 0 4240 0 5 4 0 0 5
1000 712
1000 576
1083 576
1083 539
1105 539
3 3 3 0 0 4224 0 6 5 0 0 4
743 805
936 805
936 721
954 721
3 2 4 0 0 4224 0 7 5 0 0 2
744 712
955 712
3 1 5 0 0 4224 0 8 5 0 0 4
743 613
941 613
941 703
954 703
0 2 6 0 0 4096 0 0 6 10 0 3
584 604
584 814
698 814
0 1 7 0 0 4096 0 0 6 8 0 3
638 703
638 796
698 796
0 2 8 0 0 4096 0 0 7 9 0 3
669 622
669 721
699 721
0 1 7 0 0 8192 0 0 7 17 0 3
294 327
294 703
699 703
0 2 8 0 0 0 0 0 8 20 0 3
654 529
654 622
698 622
0 1 6 0 0 8192 0 0 8 21 0 3
444 511
444 604
698 604
3 1 9 0 0 4224 0 9 12 0 0 5
1059 372
1085 372
1085 382
1097 382
1097 374
3 2 10 0 0 8320 0 10 9 0 0 4
986 468
1005 468
1005 381
1013 381
3 1 11 0 0 8320 0 11 9 0 0 4
967 265
1005 265
1005 363
1013 363
0 2 12 0 0 8320 0 0 10 30 0 5
180 108
180 552
917 552
917 477
941 477
3 1 13 0 0 4224 0 13 10 0 0 2
865 459
941 459
3 1 14 0 0 4224 0 16 11 0 0 2
863 256
922 256
2 2 7 0 0 8320 0 21 11 0 0 5
202 159
202 327
886 327
886 274
922 274
3 2 15 0 0 4224 0 14 13 0 0 4
745 520
811 520
811 468
819 468
3 1 16 0 0 4224 0 15 13 0 0 4
744 422
811 422
811 450
819 450
0 2 8 0 0 4224 0 0 14 28 0 3
472 225
472 529
700 529
0 1 6 0 0 8192 0 0 14 27 0 3
331 297
331 511
700 511
0 2 17 0 0 8192 0 0 15 26 0 3
514 315
514 431
699 431
0 1 18 0 0 8192 0 0 15 29 0 3
371 207
371 413
699 413
3 2 19 0 0 4224 0 17 16 0 0 4
740 306
809 306
809 265
817 265
3 1 20 0 0 4224 0 18 16 0 0 4
735 216
809 216
809 247
817 247
2 2 17 0 0 8320 0 19 17 0 0 3
494 152
494 315
695 315
0 1 6 0 0 8320 0 0 17 32 0 3
301 106
301 297
695 297
0 2 8 0 0 0 0 0 18 31 0 3
452 103
452 225
690 225
2 1 18 0 0 8320 0 20 18 0 0 3
345 154
345 207
690 207
1 1 12 0 0 0 0 3 21 0 0 3
177 108
202 108
202 123
1 1 8 0 0 0 0 1 19 0 0 3
435 103
494 103
494 116
1 1 6 0 0 0 0 2 20 0 0 3
293 106
345 106
345 118
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
761 91 934 115
771 99 923 115
19 Borrow = BC+A'C+A'B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
933 63 986 87
943 71 975 87
4 +BC)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
760 62 957 86
770 70 946 86
22 D = A'(B'C+BC')+A(B'C'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
756 27 913 51
766 35 902 51
17 Logic Equatiions:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
473 891 654 915
483 899 643 915
20 Fig: Full Subtractor
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1095 447 1164 471
1105 455 1153 471
6 Borrow
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1087 273 1116 297
1097 281 1105 297
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
405 32 434 56
415 40 423 56
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
279 34 308 58
289 42 297 58
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
126 39 155 63
136 47 144 63
1 A
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
