CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 77 191 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44092.5 0
0
13 Logic Switch~
5 79 131 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44092.5 0
0
14 Logic Display~
6 761 308 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3124 0 0
2
44092.5 0
0
9 2-In NOR~
219 501 331 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3421 0 0
2
44092.5 0
0
5 4049~
219 498 164 0 2 22
0 6 5
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
8157 0 0
2
44092.5 0
0
14 Logic Display~
6 764 147 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
44092.5 0
0
8 2-In OR~
219 252 168 0 3 22
0 4 3 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8901 0 0
2
44092.5 0
0
7
3 1 2 0 0 4224 0 4 3 0 0 3
540 331
761 331
761 326
0 2 3 0 0 8320 0 0 4 6 0 3
207 191
207 340
488 340
0 1 4 0 0 8320 0 0 4 7 0 3
188 131
188 322
488 322
2 1 5 0 0 4224 0 5 6 0 0 5
519 164
752 164
752 173
764 173
764 165
3 1 6 0 0 4224 0 7 5 0 0 4
285 168
475 168
475 164
483 164
1 2 3 0 0 128 0 1 7 0 0 4
89 191
231 191
231 177
239 177
1 1 4 0 0 128 0 2 7 0 0 4
91 131
231 131
231 159
239 159
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
466 417 591 441
476 425 580 441
13 Fig: NOR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
608 292 677 316
618 300 666 316
6 (A+B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
812 291 985 315
822 299 974 315
19 Using NOR Gate Chip
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
976 131 1037 155
986 139 1026 155
5 Gates
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
808 130 989 154
818 138 978 154
20 NOR Gate Using Basic
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
602 123 671 147
612 131 660 147
6 (A+B)'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
343 128 388 152
353 136 377 152
3 A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
68 197 97 221
78 205 86 221
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
67 74 96 98
77 82 85 98
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
