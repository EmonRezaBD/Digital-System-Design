CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
320 0 30 100 10
176 80 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 541 100 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89953e-315 0
0
13 Logic Switch~
5 391 98 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89953e-315 0
0
14 Logic Display~
6 1171 417 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.89953e-315 0
0
9 2-In AND~
219 816 435 0 3 22
0 4 3 2
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3421 0 0
2
5.89953e-315 0
0
14 Logic Display~
6 1150 203 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89953e-315 0
0
8 2-In OR~
219 976 229 0 3 22
0 7 6 5
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
5.89953e-315 0
0
9 Inverter~
13 597 139 0 2 22
0 3 8
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
8901 0 0
2
5.89953e-315 0
0
9 Inverter~
13 435 138 0 2 22
0 9 4
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7361 0 0
2
5.89953e-315 0
0
9 2-In AND~
219 814 308 0 3 22
0 9 8 6
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4747 0 0
2
5.89953e-315 0
0
9 2-In AND~
219 811 156 0 3 22
0 4 3 7
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
5.89953e-315 0
0
12
3 1 2 0 0 4224 0 4 3 0 0 2
837 435
1171 435
0 2 3 0 0 4224 0 0 4 10 0 3
564 100
564 444
792 444
0 1 4 0 0 8192 0 0 4 11 0 3
464 157
464 426
792 426
3 1 5 0 0 4224 0 6 5 0 0 3
1009 229
1150 229
1150 221
3 2 6 0 0 4224 0 9 6 0 0 4
835 308
955 308
955 238
963 238
3 1 7 0 0 4224 0 10 6 0 0 4
832 156
955 156
955 220
963 220
0 1 3 0 0 0 0 0 7 10 0 2
600 100
600 121
2 2 8 0 0 8320 0 7 9 0 0 3
600 157
600 317
790 317
0 1 9 0 0 8320 0 0 9 12 0 3
410 98
410 299
790 299
1 2 3 0 0 0 0 1 10 0 0 4
553 100
774 100
774 165
787 165
2 1 4 0 0 8320 0 8 10 0 0 5
438 156
438 157
779 157
779 147
787 147
1 1 9 0 0 0 0 2 8 0 0 3
403 98
438 98
438 120
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
969 76 1086 100
979 84 1075 100
12 Borrow = A'B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1074 52 1151 76
1084 60 1140 76
7 A'B+AB'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
969 53 1086 77
979 61 1075 77
12 Difference =
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
958 22 1107 46
968 30 1096 46
16 Logic Equations:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
380 32 409 56
390 40 398 56
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
537 30 566 54
547 38 555 54
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1158 353 1227 377
1168 361 1216 377
6 Borrow
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1144 143 1245 167
1154 151 1234 167
10 Difference
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
568 540 621 564
578 548 610 564
4 Fig:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
619 540 760 564
629 548 749 564
15 Half Subtractor
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
