CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 48 151 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44082.4 0
0
13 Logic Switch~
5 266 145 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44082.4 0
0
13 Logic Switch~
5 183 148 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44082.4 0
0
13 Logic Switch~
5 111 150 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
44082.4 0
0
14 Logic Display~
6 601 434 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
44082.4 0
0
14 Logic Display~
6 599 296 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
44082.4 0
0
14 Logic Display~
6 599 170 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
44082.4 0
0
8 4-In OR~
219 482 454 0 5 22
0 8 7 6 5 2
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
7361 0 0
2
44082.4 0
0
8 3-In OR~
219 474 321 0 4 22
0 8 7 6 3
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
4747 0 0
2
44082.4 0
0
8 2-In OR~
219 473 198 0 3 22
0 8 7 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
44082.4 0
0
12
5 1 2 0 0 4224 0 8 5 0 0 5
515 454
589 454
589 460
601 460
601 452
4 1 3 0 0 4224 0 9 6 0 0 3
507 321
599 321
599 314
3 1 4 0 0 4224 0 10 7 0 0 3
506 198
599 198
599 188
4 1 5 0 0 4224 0 8 1 0 0 6
465 468
79 468
79 152
63 152
63 151
60 151
0 3 6 0 0 8192 0 0 8 10 0 3
277 330
277 459
465 459
0 2 7 0 0 4112 0 0 8 8 0 3
363 321
363 450
465 450
0 1 8 0 0 4096 0 0 8 9 0 3
427 312
427 441
465 441
0 2 7 0 0 8192 0 0 9 11 0 3
310 207
310 321
462 321
0 1 8 0 0 0 0 0 9 12 0 3
409 170
409 312
461 312
1 3 6 0 0 12416 0 4 9 0 0 4
123 150
144 150
144 330
461 330
1 2 7 0 0 12416 0 3 10 0 0 4
195 148
208 148
208 207
460 207
1 1 8 0 0 8320 0 2 10 0 0 4
278 145
278 170
460 170
460 189
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
667 414 744 438
677 422 733 438
7 4-In OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
668 299 745 323
678 307 734 323
7 3-In OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
664 173 741 197
674 181 730 197
7 2-In OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
250 75 279 99
260 83 268 99
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
174 78 203 102
184 86 192 102
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
107 80 136 104
117 88 125 104
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
40 81 69 105
50 89 58 105
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
516 75 593 99
526 83 582 99
7 OR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
503 38 612 62
513 46 601 62
11 Basic Gates
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
